Library ieee;
Use ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

Entity lab6 Is
	port ( Clkin : in std_logic;
			clkout : out std_logic);
End lab6;


ARCHITECTURE Bee OF lab6 is
signal count : unsigned(19 downto 0) := "00000000000000000000";
begin 
Process (Clkin)
BEGIN 
	If (Clkin'event and Clkin ='1') then 
		count <= count+1;
	end if;
	end process;
	 clkout <= count(19);
END Bee;
